module comb_assign(
    input clk,
    input rst,
    input a,
    output b
);

    assign b = a;

endmodule
